** Profile: "SCHEMATIC1-tasi"  [ C:\Users\Ilias\Desktop\spice\ergasia-PSpiceFiles\SCHEMATIC1\tasi.sim ] 

** Creating circuit file "tasi.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Ilias\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 0.002 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
